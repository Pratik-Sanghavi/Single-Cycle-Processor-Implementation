// STAGE 2: INSTRUCTION DECODE UNIT:
// Will generate the Data signals to be delivered to ALU
// Houses the register which may be modified in the write back stage
// Control signals in this unit include reset,RegWrite, Imm_Sel, Write_Data
 
module Instruction_Decode(clk, reset, Instruction_Code, RegWrite, Imm_Sel, Write_Data, Read_Data_1, Read_Data_2, Gen_Imm_Data);

//Declaration of inputs of the decode unit
input clk;
input reset;
input [31:0]Instruction_Code; // from the Instruction Fetch Unit; will be connected later
input RegWrite; //will be generated by the control unit
input Imm_Sel; //from main control unit; facilitates mapping of input immediate data bits as per instruction format to appropriate loaction for further operations
input [31:0] Write_Data; //will be generated during the write back stage

// Declaration of outputs of the decode unit
output [31:0] Read_Data_1;
output [31:0] Read_Data_2;
output [31:0] Gen_Imm_Data;

// internal connections in the instruction decode segment
wire [4:0]Read_Register_1;
wire [4:0]Read_Register_2;
wire [4:0]Write_Register;

//Assign appropriate bits as per the rs1, rs2 and rd fields to the intermediary wires
assign Read_Register_1=Instruction_Code[20:16];
assign Read_Register_2=Instruction_Code[15:11];
assign Write_Register=Instruction_Code[25:21];

// Instantiate the Register file
Register_file RF(Read_Register_1, Read_Register_2, Write_Register, Write_Data, RegWrite, clk, reset, Read_Data_1, Read_Data_2);

// Instantiate the immediate generation unit
Immediate_Generate IG(Instruction_Code[20:0], Imm_Sel, Gen_Imm_Data); //Generates the sign extended immediate data as per instruction type

endmodule